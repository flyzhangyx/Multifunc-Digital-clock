library verilog;
use verilog.vl_types.all;
entity cntall_vlg_vec_tst is
end cntall_vlg_vec_tst;
