library verilog;
use verilog.vl_types.all;
entity cnt6_vlg_vec_tst is
end cnt6_vlg_vec_tst;
