library verilog;
use verilog.vl_types.all;
entity Do_vlg_sample_tst is
    port(
        clik            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Do_vlg_sample_tst;
