library verilog;
use verilog.vl_types.all;
entity switchlll_vlg_vec_tst is
end switchlll_vlg_vec_tst;
