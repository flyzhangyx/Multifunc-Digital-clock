library verilog;
use verilog.vl_types.all;
entity boom_vlg_vec_tst is
end boom_vlg_vec_tst;
