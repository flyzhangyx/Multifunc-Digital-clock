library verilog;
use verilog.vl_types.all;
entity cnt8_vlg_vec_tst is
end cnt8_vlg_vec_tst;
