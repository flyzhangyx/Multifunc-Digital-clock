library verilog;
use verilog.vl_types.all;
entity m200_vlg_vec_tst is
end m200_vlg_vec_tst;
