library verilog;
use verilog.vl_types.all;
entity dig_select_vlg_vec_tst is
end dig_select_vlg_vec_tst;
