library verilog;
use verilog.vl_types.all;
entity switchlll_vlg_check_tst is
    port(
        key_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end switchlll_vlg_check_tst;
