library verilog;
use verilog.vl_types.all;
entity Do_vlg_vec_tst is
end Do_vlg_vec_tst;
