library verilog;
use verilog.vl_types.all;
entity m200_vlg_check_tst is
    port(
        carry           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end m200_vlg_check_tst;
