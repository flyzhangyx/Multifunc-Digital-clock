library verilog;
use verilog.vl_types.all;
entity m100 is
    port(
        co              : out    vl_logic;
        clk             : in     vl_logic
    );
end m100;
