library verilog;
use verilog.vl_types.all;
entity timedelay_vlg_vec_tst is
end timedelay_vlg_vec_tst;
