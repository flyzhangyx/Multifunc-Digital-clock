library verilog;
use verilog.vl_types.all;
entity Do_vlg_check_tst is
    port(
        clik_250hz      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Do_vlg_check_tst;
