library verilog;
use verilog.vl_types.all;
entity chooseseg_vlg_vec_tst is
end chooseseg_vlg_vec_tst;
