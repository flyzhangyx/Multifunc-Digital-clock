library verilog;
use verilog.vl_types.all;
entity music_vlg_vec_tst is
end music_vlg_vec_tst;
