library verilog;
use verilog.vl_types.all;
entity decoder_vlg_vec_tst is
end decoder_vlg_vec_tst;
