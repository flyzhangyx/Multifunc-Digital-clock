library verilog;
use verilog.vl_types.all;
entity music_vlg_check_tst is
    port(
        music           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end music_vlg_check_tst;
