library verilog;
use verilog.vl_types.all;
entity boom_vlg_check_tst is
    port(
        delay           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end boom_vlg_check_tst;
