library verilog;
use verilog.vl_types.all;
entity choose_vlg_vec_tst is
end choose_vlg_vec_tst;
