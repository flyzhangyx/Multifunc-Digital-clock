library verilog;
use verilog.vl_types.all;
entity choose_vlg_check_tst is
    port(
        outputdig       : in     vl_logic_vector(5 downto 0);
        sampler_rx      : in     vl_logic
    );
end choose_vlg_check_tst;
